interface dff_if;
  logic clk;  // clock signal
  logic rst;  // Reset signal
  logic din;  // Data input
  logic dout; // Data output
endinterface
